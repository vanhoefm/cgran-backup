// -*- verilog -*-
//
//  Sensing and Processing Across Networks (SPAN) Lab.
//  University of Utah, UT-84112
//  802.11b receiver v1.0
//  Author: Mohammad H. Firooz   mhfirooz@yahoo.com
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation; either version 2 of the License, or
//  (at your option) any later version.
//
//  This program is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this program; if not, write to the Free Software
//  Foundation, Inc., 51 Franklin Street, Boston, MA  02110-1301  USA
//


module ComplexAbs(datai, dataq, absval);
input [15:0] datai, dataq;
output [32:0] absval;

wire [31:0] datai2, dataq2;
power2 power2i(
	.dataa(datai),
	.result(datai2));

power2 power2q(
	.dataa(dataq),
	.result(dataq2));
	
padd52 adder(
	.data0x(dataq2),
	.data1x(datai2),
	.result(absval));


endmodule

// megafunction wizard: %LPM_ABS%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_abs 

// ============================================================
// File Name: singleABS.v
// Megafunction Name(s):
// 			lpm_abs
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Build 175 11/20/2007 SP 1 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module singleABS (
	data,
	result);

	input	[25:0]  data;
	output	[25:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone"
// Retrieval info: PRIVATE: OptionalOverflowOutput NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: nBit NUMERIC "26"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_ABS"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "26"
// Retrieval info: USED_PORT: data 0 0 26 0 INPUT NODEFVAL data[25..0]
// Retrieval info: USED_PORT: result 0 0 26 0 OUTPUT NODEFVAL result[25..0]
// Retrieval info: CONNECT: @data 0 0 26 0 data 0 0 26 0
// Retrieval info: CONNECT: result 0 0 26 0 @result 0 0 26 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL singleABS_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
